module bcd7seg(
  input  [3:0] b,
  output reg [6:0] h
);

always @(*) begin
  case (b)
    4'b0000: h = 7'b0000001; // 0
    4'b0001: h = 7'b1001111; // 1
    4'b0010: h = 7'b0010010; // 2
    4'b0011: h = 7'b0000110; // 3
    4'b0100: h = 7'b1001100; // 4
    4'b0101: h = 7'b0100100; // 5
    4'b0110: h = 7'b0100000; // 6
    4'b0111: h = 7'b0001111; // 7
    4'b1000: h = 7'b0000000; // 8
    4'b1001: h = 7'b0000100; // 9
    default: h = 7'b0000000; // off
  endcase
end
endmodule

